// look in pins.pcf for all the pin names on the TinyFPGA BX board

module hera (
  input [15:0] opcode,
  output [15:0]

  );

endmodule // hera



module top (
    input CLK,    // 16MHz clock
    output LED,   // User/boot LED next to power LED



);


endmodule
